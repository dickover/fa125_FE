--  C:\USERS\DICKOVER\DOCUMENTS\...\FT_PROCESSM_CDC_FDC.vhd
--  VHDL code created by Xilinx's StateCAD 10.1
--  Fri Mar 11 13:02:31 2016

--  This VHDL code (for use with Xilinx XST) was generated using: 
--  enumerated state assignment with structured code format.
--  Minimization is enabled,  implied else is enabled, 
--  and outputs are speed optimized.

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SHELL_FT_PROCESSM_CDC_FDC IS
	PORT (CLK,FT_ABOVE_TH,FT_DONE,GO,INIT_PED_CALC_DN,LOC_PED_CALC_DN,MODE0,
		MODE1,MODE2,NO_EVENT,PEAK_WRITE_DONE,PTW_DONE,RESET_N,wait_PG_done,WE_DONE: 
		IN std_logic;
		CLR_INIT_PED_CNT,CLR_LOC_PED_CNT,CLR_PTW_DONE,DEC_PEAK_CNT,FT_GO,
			HOST_BLOCK_INC,IDLE,LatchNoEvenClr,NoEventLatch,NOT_VALID_2,PINIT_CALC_EN,
			PLOCAL_CALC_EN,PR_FIFO_WR_EN,PR_FIFO_WR_EN_TR,PTW_CNT_CLR,RAW_PTW_PTR_EN,
			RD_PTW_PTR_EN_5,RT_PTW_PTR,RT_PTW_PTR_2,RT_PTW_PTR_PLOC,SAVE_PTW_PTR,
			SAVE_PTW_PTR_FT,SEL_CDC_FT_WD_1,SEL_CDC_FT_WD_2,SEL_FDC_AMP_WD_1,
			SEL_FDC_AMP_WD_2,SEL_FDC_SUM_WD_1,SEL_FDC_SUM_WD_2,SEL_RAW_SAMPLE_2,SEL_RS_1,
			SEL_RS_2,SEL_WIN_RAW_WD_1 : OUT std_logic);
END;

ARCHITECTURE BEHAVIOR OF SHELL_FT_PROCESSM_CDC_FDC IS
	TYPE type_sreg IS (ADJUSTCNT,Choose_mode,CruisePTWBuf,Main_IDLE,MAIN_WAIT1,
		MAIN_WAIT2,MAIN_WAIT3,STATE1,STATE23);
	SIGNAL sreg, next_sreg : type_sreg;
	TYPE type_sreg1 IS (MODE_IDLE,Pulse_Data,PULSE_DATA_END,STATE0,STATE3,STATE4
		,STATE5,STATE6,STATE7,STATE8,STATE9,STATE10,STATE11,STATE12,STATE13,STATE15,
		STATE19,STATE21,STATE22,STATE24,STATE25,STATE26,STATE27,STATE28,STATE30,
		STATE31,STATE32,STATE33,STATE35,STATE36,STATE37,STATE38,STATE41,STATE42,
		STATE43,STATE44,STATE45,STATE46,STATE47,STATE48,STATE49,STATE50,STATE51,
		STATE53,STATE54,STATE55,STATE56,STATE57,STATE58,STATE59,STATE60,STATE61,
		STATE62,STATE63,STATE64,STATE65,STATE66,STATE69,STATE70,STATE71,STATE72,
		STATE73,STATE74,STATE75,STATE77,STATE78,STATE79,STATE80,STATE81,STATE82);
	SIGNAL sreg1, next_sreg1 : type_sreg1;
	TYPE type_sreg2 IS (Cruise_Done_FT,Cruise_Mode,CRUISEBUFFER_FT,CruiseIdle,
		FT_HAVE_DATA,FT_NODATA,PINIT_cruise_DLY,PINT_CALC,PLOCAL_CALC,RestorePTR_FT,
		STATE2,STATE14,STATE16,STATE17,STATE18,STATE20,STATE29,STATE39,STATE40,
		STATE52,STATE67);
	SIGNAL sreg2, next_sreg2 : type_sreg2;
	SIGNAL next_CLR_INIT_PED_CNT,next_CLR_LOC_PED_CNT,next_CLR_PTW_DONE,
		next_CruiseDone,next_CruiseON,next_DEC_PEAK_CNT,next_FT_GO,
		next_HOST_BLOCK_INC,next_IDLE,next_LatchNoEvenClr,next_MODE_DONE,next_MODE_GO
		,next_NoEventLatch,next_NOT_VALID_2,next_PINIT_CALC_EN,next_PLOCAL_CALC_EN,
		next_PR_FIFO_WR_EN,next_PR_FIFO_WR_EN_TR,next_PTW_CNT_CLR,next_RAW_PTW_PTR_EN
		,next_RD_PTW_PTR_EN_5,next_RT_PTW_PTR,next_RT_PTW_PTR_2,next_RT_PTW_PTR_PLOC,
		next_SAVE_PTW_PTR,next_SAVE_PTW_PTR_FT,next_SEL_CDC_FT_WD_1,
		next_SEL_CDC_FT_WD_2,next_SEL_FDC_AMP_WD_1,next_SEL_FDC_AMP_WD_2,
		next_SEL_FDC_SUM_WD_1,next_SEL_FDC_SUM_WD_2,next_SEL_RAW_SAMPLE_2,
		next_SEL_RS_1,next_SEL_RS_2,next_SEL_WIN_RAW_WD_1 : std_logic;

	SIGNAL CruiseDone,CruiseON,MODE_DONE,MODE_GO: std_logic;
BEGIN
	PROCESS (CLK, next_sreg, next_CLR_PTW_DONE, next_CruiseON, 
		next_HOST_BLOCK_INC, next_IDLE, next_LatchNoEvenClr, next_MODE_GO, 
		next_PR_FIFO_WR_EN_TR, next_SAVE_PTW_PTR)
	BEGIN
		IF CLK='1' AND CLK'event THEN
			sreg <= next_sreg;
			CLR_PTW_DONE <= next_CLR_PTW_DONE;
			CruiseON <= next_CruiseON;
			HOST_BLOCK_INC <= next_HOST_BLOCK_INC;
			IDLE <= next_IDLE;
			LatchNoEvenClr <= next_LatchNoEvenClr;
			MODE_GO <= next_MODE_GO;
			PR_FIFO_WR_EN_TR <= next_PR_FIFO_WR_EN_TR;
			SAVE_PTW_PTR <= next_SAVE_PTW_PTR;
		END IF;
	END PROCESS;

	PROCESS (CLK, next_sreg1, next_DEC_PEAK_CNT, next_FT_GO, next_MODE_DONE, 
		next_NOT_VALID_2, next_PR_FIFO_WR_EN, next_RAW_PTW_PTR_EN, next_RT_PTW_PTR_2,
		 next_SEL_CDC_FT_WD_1, next_SEL_CDC_FT_WD_2, next_SEL_FDC_AMP_WD_1, 
		next_SEL_FDC_AMP_WD_2, next_SEL_FDC_SUM_WD_1, next_SEL_FDC_SUM_WD_2, 
		next_SEL_RAW_SAMPLE_2, next_SEL_RS_1, next_SEL_RS_2, next_SEL_WIN_RAW_WD_1)
	BEGIN
		IF CLK='1' AND CLK'event THEN
			sreg1 <= next_sreg1;
			DEC_PEAK_CNT <= next_DEC_PEAK_CNT;
			FT_GO <= next_FT_GO;
			MODE_DONE <= next_MODE_DONE;
			NOT_VALID_2 <= next_NOT_VALID_2;
			PR_FIFO_WR_EN <= next_PR_FIFO_WR_EN;
			RAW_PTW_PTR_EN <= next_RAW_PTW_PTR_EN;
			RT_PTW_PTR_2 <= next_RT_PTW_PTR_2;
			SEL_CDC_FT_WD_1 <= next_SEL_CDC_FT_WD_1;
			SEL_CDC_FT_WD_2 <= next_SEL_CDC_FT_WD_2;
			SEL_FDC_AMP_WD_1 <= next_SEL_FDC_AMP_WD_1;
			SEL_FDC_AMP_WD_2 <= next_SEL_FDC_AMP_WD_2;
			SEL_FDC_SUM_WD_1 <= next_SEL_FDC_SUM_WD_1;
			SEL_FDC_SUM_WD_2 <= next_SEL_FDC_SUM_WD_2;
			SEL_RAW_SAMPLE_2 <= next_SEL_RAW_SAMPLE_2;
			SEL_RS_1 <= next_SEL_RS_1;
			SEL_RS_2 <= next_SEL_RS_2;
			SEL_WIN_RAW_WD_1 <= next_SEL_WIN_RAW_WD_1;
		END IF;
	END PROCESS;

	PROCESS (CLK, next_sreg2, next_CLR_INIT_PED_CNT, next_CLR_LOC_PED_CNT, 
		next_CruiseDone, next_NoEventLatch, next_PINIT_CALC_EN, next_PLOCAL_CALC_EN, 
		next_PTW_CNT_CLR, next_RD_PTW_PTR_EN_5, next_RT_PTW_PTR, next_RT_PTW_PTR_PLOC
		, next_SAVE_PTW_PTR_FT)
	BEGIN
		IF CLK='1' AND CLK'event THEN
			sreg2 <= next_sreg2;
			CLR_INIT_PED_CNT <= next_CLR_INIT_PED_CNT;
			CLR_LOC_PED_CNT <= next_CLR_LOC_PED_CNT;
			CruiseDone <= next_CruiseDone;
			NoEventLatch <= next_NoEventLatch;
			PINIT_CALC_EN <= next_PINIT_CALC_EN;
			PLOCAL_CALC_EN <= next_PLOCAL_CALC_EN;
			PTW_CNT_CLR <= next_PTW_CNT_CLR;
			RD_PTW_PTR_EN_5 <= next_RD_PTW_PTR_EN_5;
			RT_PTW_PTR <= next_RT_PTW_PTR;
			RT_PTW_PTR_PLOC <= next_RT_PTW_PTR_PLOC;
			SAVE_PTW_PTR_FT <= next_SAVE_PTW_PTR_FT;
		END IF;
	END PROCESS;

	PROCESS (sreg,sreg1,sreg2,CruiseDone,CruiseON,FT_ABOVE_TH,FT_DONE,GO,
		INIT_PED_CALC_DN,LOC_PED_CALC_DN,MODE0,MODE1,MODE2,MODE_DONE,MODE_GO,NO_EVENT
		,PEAK_WRITE_DONE,PTW_DONE,RESET_N,wait_PG_done,WE_DONE)
	BEGIN
		next_CLR_INIT_PED_CNT <= '0'; next_CLR_LOC_PED_CNT <= '0'; 
			next_CLR_PTW_DONE <= '0'; next_CruiseDone <= '0'; next_CruiseON <= '0'; 
			next_DEC_PEAK_CNT <= '0'; next_FT_GO <= '0'; next_HOST_BLOCK_INC <= '0'; 
			next_IDLE <= '0'; next_LatchNoEvenClr <= '0'; next_MODE_DONE <= '0'; 
			next_MODE_GO <= '0'; next_NoEventLatch <= '0'; next_NOT_VALID_2 <= '0'; 
			next_PINIT_CALC_EN <= '0'; next_PLOCAL_CALC_EN <= '0'; next_PR_FIFO_WR_EN <= 
			'0'; next_PR_FIFO_WR_EN_TR <= '0'; next_PTW_CNT_CLR <= '0'; 
			next_RAW_PTW_PTR_EN <= '0'; next_RD_PTW_PTR_EN_5 <= '0'; next_RT_PTW_PTR <= 
			'0'; next_RT_PTW_PTR_2 <= '0'; next_RT_PTW_PTR_PLOC <= '0'; next_SAVE_PTW_PTR
			 <= '0'; next_SAVE_PTW_PTR_FT <= '0'; next_SEL_CDC_FT_WD_1 <= '0'; 
			next_SEL_CDC_FT_WD_2 <= '0'; next_SEL_FDC_AMP_WD_1 <= '0'; 
			next_SEL_FDC_AMP_WD_2 <= '0'; next_SEL_FDC_SUM_WD_1 <= '0'; 
			next_SEL_FDC_SUM_WD_2 <= '0'; next_SEL_RAW_SAMPLE_2 <= '0'; next_SEL_RS_1 <= 
			'0'; next_SEL_RS_2 <= '0'; next_SEL_WIN_RAW_WD_1 <= '0'; 

		next_sreg<=ADJUSTCNT;
		next_sreg1<=MODE_IDLE;
		next_sreg2<=Cruise_Done_FT;

		IF ( RESET_N='0' ) THEN
			next_sreg<=Main_IDLE;
			next_CruiseON<='0';
			next_HOST_BLOCK_INC<='0';
			next_LatchNoEvenClr<='0';
			next_MODE_GO<='0';
			next_PR_FIFO_WR_EN_TR<='0';
			next_CLR_PTW_DONE<='1';
			next_SAVE_PTW_PTR<='1';
			next_IDLE<='1';
		ELSE
			CASE sreg IS
				WHEN ADJUSTCNT =>
					next_sreg<=MAIN_WAIT1;
					next_CLR_PTW_DONE<='0';
					next_CruiseON<='0';
					next_HOST_BLOCK_INC<='0';
					next_IDLE<='0';
					next_MODE_GO<='0';
					next_PR_FIFO_WR_EN_TR<='0';
					next_SAVE_PTW_PTR<='0';
					next_LatchNoEvenClr<='1';
				WHEN Choose_mode =>
					IF ( MODE_DONE='1' ) THEN
						next_sreg<=STATE23;
						next_CLR_PTW_DONE<='0';
						next_CruiseON<='0';
						next_HOST_BLOCK_INC<='0';
						next_IDLE<='0';
						next_LatchNoEvenClr<='0';
						next_MODE_GO<='0';
						next_SAVE_PTW_PTR<='0';
						next_PR_FIFO_WR_EN_TR<='1';
					 ELSE
						next_sreg<=Choose_mode;
						next_CLR_PTW_DONE<='0';
						next_CruiseON<='0';
						next_HOST_BLOCK_INC<='0';
						next_IDLE<='0';
						next_LatchNoEvenClr<='0';
						next_PR_FIFO_WR_EN_TR<='0';
						next_SAVE_PTW_PTR<='0';
						next_MODE_GO<='1';
					END IF;
				WHEN CruisePTWBuf =>
					IF ( CruiseDone='1' ) THEN
						next_sreg<=STATE1;
						next_CLR_PTW_DONE<='0';
						next_CruiseON<='0';
						next_HOST_BLOCK_INC<='0';
						next_IDLE<='0';
						next_LatchNoEvenClr<='0';
						next_MODE_GO<='0';
						next_PR_FIFO_WR_EN_TR<='0';
						next_SAVE_PTW_PTR<='0';
					 ELSE
						next_sreg<=CruisePTWBuf;
						next_CLR_PTW_DONE<='0';
						next_HOST_BLOCK_INC<='0';
						next_IDLE<='0';
						next_LatchNoEvenClr<='0';
						next_MODE_GO<='0';
						next_PR_FIFO_WR_EN_TR<='0';
						next_SAVE_PTW_PTR<='0';
						next_CruiseON<='1';
					END IF;
				WHEN Main_IDLE =>
					IF ( GO='1' ) THEN
						next_sreg<=CruisePTWBuf;
						next_CLR_PTW_DONE<='0';
						next_HOST_BLOCK_INC<='0';
						next_IDLE<='0';
						next_LatchNoEvenClr<='0';
						next_MODE_GO<='0';
						next_PR_FIFO_WR_EN_TR<='0';
						next_SAVE_PTW_PTR<='0';
						next_CruiseON<='1';
					 ELSE
						next_sreg<=Main_IDLE;
						next_CruiseON<='0';
						next_HOST_BLOCK_INC<='0';
						next_LatchNoEvenClr<='0';
						next_MODE_GO<='0';
						next_PR_FIFO_WR_EN_TR<='0';
						next_CLR_PTW_DONE<='1';
						next_SAVE_PTW_PTR<='1';
						next_IDLE<='1';
					END IF;
				WHEN MAIN_WAIT1 =>
					next_sreg<=MAIN_WAIT2;
					next_CLR_PTW_DONE<='0';
					next_CruiseON<='0';
					next_HOST_BLOCK_INC<='0';
					next_IDLE<='0';
					next_LatchNoEvenClr<='0';
					next_MODE_GO<='0';
					next_PR_FIFO_WR_EN_TR<='0';
					next_SAVE_PTW_PTR<='0';
				WHEN MAIN_WAIT2 =>
					next_sreg<=MAIN_WAIT3;
					next_CLR_PTW_DONE<='0';
					next_CruiseON<='0';
					next_HOST_BLOCK_INC<='0';
					next_LatchNoEvenClr<='0';
					next_MODE_GO<='0';
					next_PR_FIFO_WR_EN_TR<='0';
					next_SAVE_PTW_PTR<='0';
					next_IDLE<='1';
				WHEN MAIN_WAIT3 =>
					next_sreg<=Main_IDLE;
					next_CruiseON<='0';
					next_HOST_BLOCK_INC<='0';
					next_LatchNoEvenClr<='0';
					next_MODE_GO<='0';
					next_PR_FIFO_WR_EN_TR<='0';
					next_CLR_PTW_DONE<='1';
					next_SAVE_PTW_PTR<='1';
					next_IDLE<='1';
				WHEN STATE1 =>
					IF ( NO_EVENT='0' ) THEN
						next_sreg<=Choose_mode;
						next_CLR_PTW_DONE<='0';
						next_CruiseON<='0';
						next_HOST_BLOCK_INC<='0';
						next_IDLE<='0';
						next_LatchNoEvenClr<='0';
						next_PR_FIFO_WR_EN_TR<='0';
						next_SAVE_PTW_PTR<='0';
						next_MODE_GO<='1';
					END IF;
					IF ( NO_EVENT='1' ) THEN
						next_sreg<=STATE23;
						next_CLR_PTW_DONE<='0';
						next_CruiseON<='0';
						next_HOST_BLOCK_INC<='0';
						next_IDLE<='0';
						next_LatchNoEvenClr<='0';
						next_MODE_GO<='0';
						next_SAVE_PTW_PTR<='0';
						next_PR_FIFO_WR_EN_TR<='1';
					END IF;
				WHEN STATE23 =>
					next_sreg<=ADJUSTCNT;
					next_CLR_PTW_DONE<='0';
					next_CruiseON<='0';
					next_IDLE<='0';
					next_LatchNoEvenClr<='0';
					next_MODE_GO<='0';
					next_PR_FIFO_WR_EN_TR<='0';
					next_SAVE_PTW_PTR<='0';
					next_HOST_BLOCK_INC<='1';
				WHEN OTHERS =>
			END CASE;
		END IF;

		IF ( RESET_N='0' ) THEN
			next_sreg1<=MODE_IDLE;
			next_DEC_PEAK_CNT<='0';
			next_FT_GO<='0';
			next_MODE_DONE<='0';
			next_NOT_VALID_2<='0';
			next_PR_FIFO_WR_EN<='0';
			next_RAW_PTW_PTR_EN<='0';
			next_RT_PTW_PTR_2<='0';
			next_SEL_CDC_FT_WD_1<='0';
			next_SEL_CDC_FT_WD_2<='0';
			next_SEL_FDC_AMP_WD_1<='0';
			next_SEL_FDC_AMP_WD_2<='0';
			next_SEL_FDC_SUM_WD_1<='0';
			next_SEL_FDC_SUM_WD_2<='0';
			next_SEL_RAW_SAMPLE_2<='0';
			next_SEL_RS_1<='0';
			next_SEL_RS_2<='0';
			next_SEL_WIN_RAW_WD_1<='0';
		ELSE
			CASE sreg1 IS
				WHEN MODE_IDLE =>
					IF ( MODE_GO='1' ) THEN
						next_sreg1<=STATE5;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
					 ELSE
						next_sreg1<=MODE_IDLE;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
					END IF;
				WHEN Pulse_Data =>
					IF ( FT_DONE='1' ) THEN
						next_sreg1<=STATE80;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_SEL_CDC_FT_WD_1<='1';
					 ELSE
						next_sreg1<=Pulse_Data;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
				WHEN PULSE_DATA_END =>
					next_sreg1<=STATE42;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE0 =>
					next_sreg1<=MODE_IDLE;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE3 =>
					IF ( PEAK_WRITE_DONE='1' ) THEN
						next_sreg1<=STATE0;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_MODE_DONE<='1';
					ELSIF ( PEAK_WRITE_DONE='0' ) THEN
						next_sreg1<=STATE55;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
					END IF;
				WHEN STATE4 =>
					next_sreg1<=STATE70;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='1';
				WHEN STATE5 =>
					IF ( MODE2='0' AND MODE1='0' ) THEN
						next_sreg1<=STATE5;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
					END IF;
					IF ( MODE0='1' AND MODE1='1' AND MODE2='1' ) THEN
						next_sreg1<=STATE54;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
					IF ( MODE0='0' AND MODE1='1' AND MODE2='1' ) THEN
						next_sreg1<=STATE12;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
					IF ( MODE0='1' AND MODE1='0' AND MODE2='1' ) THEN
						next_sreg1<=STATE46;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
					IF ( MODE1='0' AND MODE0='0' AND MODE2='1' ) THEN
						next_sreg1<=STATE35;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
					IF ( MODE2='0' AND MODE0='1' AND MODE1='1' ) THEN
						next_sreg1<=STATE30;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
					IF ( MODE2='0' AND MODE0='0' AND MODE1='1' ) THEN
						next_sreg1<=Pulse_Data;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
				WHEN STATE6 =>
					IF ( PEAK_WRITE_DONE='1' ) THEN
						next_sreg1<=STATE11;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_RT_PTW_PTR_2<='1';
						next_SEL_WIN_RAW_WD_1<='1';
					ELSIF ( PEAK_WRITE_DONE='0' ) THEN
						next_sreg1<=STATE65;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
					END IF;
				WHEN STATE7 =>
					next_sreg1<=STATE22;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE8 =>
					next_sreg1<=STATE10;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE9 =>
					next_sreg1<=STATE27;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='1';
					next_PR_FIFO_WR_EN<='1';
				WHEN STATE10 =>
					IF ( PTW_DONE='1' ) THEN
						next_sreg1<=STATE26;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_NOT_VALID_2<='1';
					ELSIF ( PTW_DONE='0' ) THEN
						next_sreg1<=STATE25;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_SEL_RS_2<='1';
						next_RAW_PTW_PTR_EN<='1';
					END IF;
				WHEN STATE11 =>
					next_sreg1<=STATE7;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='1';
					next_PR_FIFO_WR_EN<='1';
				WHEN STATE12 =>
					IF ( FT_DONE='1' ) THEN
						next_sreg1<=STATE79;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_SEL_FDC_SUM_WD_1<='1';
					 ELSE
						next_sreg1<=STATE12;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
				WHEN STATE13 =>
					next_sreg1<=STATE74;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='1';
				WHEN STATE15 =>
					next_sreg1<=STATE49;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE19 =>
					IF ( PEAK_WRITE_DONE='1' ) THEN
						next_sreg1<=STATE11;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_RT_PTW_PTR_2<='1';
						next_SEL_WIN_RAW_WD_1<='1';
					ELSIF ( PEAK_WRITE_DONE='0' ) THEN
						next_sreg1<=STATE63;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
					END IF;
				WHEN STATE21 =>
					next_sreg1<=STATE9;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='1';
				WHEN STATE22 =>
					IF ( PTW_DONE='1' ) THEN
						next_sreg1<=STATE0;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_MODE_DONE<='1';
					ELSIF ( PTW_DONE='0' ) THEN
						next_sreg1<=STATE24;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_SEL_RS_1<='1';
						next_RAW_PTW_PTR_EN<='1';
					END IF;
				WHEN STATE24 =>
					next_sreg1<=STATE8;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE25 =>
					next_sreg1<=STATE21;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE26 =>
					next_sreg1<=STATE69;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_NOT_VALID_2<='1';
				WHEN STATE27 =>
					next_sreg1<=STATE22;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE28 =>
					next_sreg1<=STATE0;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_MODE_DONE<='1';
				WHEN STATE30 =>
					IF ( FT_DONE='1' ) THEN
						next_sreg1<=STATE81;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_SEL_FDC_SUM_WD_1<='1';
					 ELSE
						next_sreg1<=STATE30;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
				WHEN STATE31 =>
					next_sreg1<=STATE71;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='1';
				WHEN STATE32 =>
					next_sreg1<=STATE43;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE33 =>
					IF ( PEAK_WRITE_DONE='1' ) THEN
						next_sreg1<=STATE0;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_MODE_DONE<='1';
					ELSIF ( PEAK_WRITE_DONE='0' ) THEN
						next_sreg1<=STATE59;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
					END IF;
				WHEN STATE35 =>
					IF ( FT_DONE='1' ) THEN
						next_sreg1<=STATE82;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_SEL_FDC_AMP_WD_1<='1';
					 ELSE
						next_sreg1<=STATE35;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
				WHEN STATE36 =>
					next_sreg1<=STATE72;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='1';
				WHEN STATE37 =>
					next_sreg1<=STATE47;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE38 =>
					IF ( PEAK_WRITE_DONE='1' ) THEN
						next_sreg1<=STATE0;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_MODE_DONE<='1';
					ELSIF ( PEAK_WRITE_DONE='0' ) THEN
						next_sreg1<=STATE57;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
					END IF;
				WHEN STATE41 =>
					next_sreg1<=STATE50;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE42 =>
					next_sreg1<=STATE3;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE43 =>
					next_sreg1<=STATE33;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE44 =>
					next_sreg1<=STATE48;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE45 =>
					next_sreg1<=STATE75;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='1';
				WHEN STATE46 =>
					IF ( FT_DONE='1' ) THEN
						next_sreg1<=STATE77;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_SEL_CDC_FT_WD_1<='1';
					 ELSE
						next_sreg1<=STATE46;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
				WHEN STATE47 =>
					next_sreg1<=STATE38;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE48 =>
					next_sreg1<=STATE6;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE49 =>
					next_sreg1<=STATE19;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE50 =>
					IF ( PEAK_WRITE_DONE='1' ) THEN
						next_sreg1<=STATE11;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_RT_PTW_PTR_2<='1';
						next_SEL_WIN_RAW_WD_1<='1';
					ELSIF ( PEAK_WRITE_DONE='0' ) THEN
						next_sreg1<=STATE61;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
					END IF;
				WHEN STATE51 =>
					next_sreg1<=STATE41;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
				WHEN STATE53 =>
					next_sreg1<=STATE73;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='1';
				WHEN STATE54 =>
					IF ( FT_DONE='1' ) THEN
						next_sreg1<=STATE78;
						next_DEC_PEAK_CNT<='0';
						next_FT_GO<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_SEL_FDC_AMP_WD_1<='1';
					 ELSE
						next_sreg1<=STATE54;
						next_DEC_PEAK_CNT<='0';
						next_MODE_DONE<='0';
						next_NOT_VALID_2<='0';
						next_PR_FIFO_WR_EN<='0';
						next_RAW_PTW_PTR_EN<='0';
						next_RT_PTW_PTR_2<='0';
						next_SEL_CDC_FT_WD_1<='0';
						next_SEL_CDC_FT_WD_2<='0';
						next_SEL_FDC_AMP_WD_1<='0';
						next_SEL_FDC_AMP_WD_2<='0';
						next_SEL_FDC_SUM_WD_1<='0';
						next_SEL_FDC_SUM_WD_2<='0';
						next_SEL_RAW_SAMPLE_2<='0';
						next_SEL_RS_1<='0';
						next_SEL_RS_2<='0';
						next_SEL_WIN_RAW_WD_1<='0';
						next_FT_GO<='1';
					END IF;
				WHEN STATE55 =>
					next_sreg1<=STATE56;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='1';
				WHEN STATE56 =>
					next_sreg1<=PULSE_DATA_END;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE57 =>
					next_sreg1<=STATE58;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='1';
				WHEN STATE58 =>
					next_sreg1<=STATE37;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE59 =>
					next_sreg1<=STATE60;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='1';
				WHEN STATE60 =>
					next_sreg1<=STATE32;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE61 =>
					next_sreg1<=STATE62;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='1';
				WHEN STATE62 =>
					next_sreg1<=STATE51;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE63 =>
					next_sreg1<=STATE64;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='1';
				WHEN STATE64 =>
					next_sreg1<=STATE15;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE65 =>
					next_sreg1<=STATE66;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_PR_FIFO_WR_EN<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='1';
				WHEN STATE66 =>
					next_sreg1<=STATE44;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE69 =>
					next_sreg1<=STATE28;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_NOT_VALID_2<='1';
				WHEN STATE70 =>
					next_sreg1<=PULSE_DATA_END;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE71 =>
					next_sreg1<=STATE32;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE72 =>
					next_sreg1<=STATE37;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE73 =>
					next_sreg1<=STATE51;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE74 =>
					next_sreg1<=STATE15;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE75 =>
					next_sreg1<=STATE44;
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='1';
					next_PR_FIFO_WR_EN<='1';
					next_DEC_PEAK_CNT<='1';
				WHEN STATE77 =>
					next_sreg1<=STATE45;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_1<='1';
					next_PR_FIFO_WR_EN<='1';
				WHEN STATE78 =>
					next_sreg1<=STATE53;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='1';
					next_PR_FIFO_WR_EN<='1';
				WHEN STATE79 =>
					next_sreg1<=STATE13;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='1';
					next_PR_FIFO_WR_EN<='1';
				WHEN STATE80 =>
					next_sreg1<=STATE4;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_CDC_FT_WD_1<='1';
					next_PR_FIFO_WR_EN<='1';
				WHEN STATE81 =>
					next_sreg1<=STATE31;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_1<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_SUM_WD_1<='1';
					next_PR_FIFO_WR_EN<='1';
				WHEN STATE82 =>
					next_sreg1<=STATE36;
					next_DEC_PEAK_CNT<='0';
					next_FT_GO<='0';
					next_MODE_DONE<='0';
					next_NOT_VALID_2<='0';
					next_RAW_PTW_PTR_EN<='0';
					next_RT_PTW_PTR_2<='0';
					next_SEL_CDC_FT_WD_1<='0';
					next_SEL_CDC_FT_WD_2<='0';
					next_SEL_FDC_AMP_WD_2<='0';
					next_SEL_FDC_SUM_WD_1<='0';
					next_SEL_FDC_SUM_WD_2<='0';
					next_SEL_RAW_SAMPLE_2<='0';
					next_SEL_RS_1<='0';
					next_SEL_RS_2<='0';
					next_SEL_WIN_RAW_WD_1<='0';
					next_SEL_FDC_AMP_WD_1<='1';
					next_PR_FIFO_WR_EN<='1';
				WHEN OTHERS =>
			END CASE;
		END IF;

		IF ( RESET_N='0' ) THEN
			next_sreg2<=CruiseIdle;
			next_CLR_INIT_PED_CNT<='0';
			next_CLR_LOC_PED_CNT<='0';
			next_CruiseDone<='0';
			next_NoEventLatch<='0';
			next_PINIT_CALC_EN<='0';
			next_PLOCAL_CALC_EN<='0';
			next_PTW_CNT_CLR<='0';
			next_RD_PTW_PTR_EN_5<='0';
			next_RT_PTW_PTR<='0';
			next_RT_PTW_PTR_PLOC<='0';
			next_SAVE_PTW_PTR_FT<='0';
		ELSE
			CASE sreg2 IS
				WHEN Cruise_Done_FT =>
					next_sreg2<=CruiseIdle;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RD_PTW_PTR_EN_5<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
				WHEN Cruise_Mode =>
					next_sreg2<=PINIT_cruise_DLY;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_RD_PTW_PTR_EN_5<='1';
				WHEN CRUISEBUFFER_FT =>
					IF ( WE_DONE='1' ) THEN
						next_sreg2<=STATE14;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RD_PTW_PTR_EN_5<='1';
					ELSIF ( FT_ABOVE_TH='1' ) THEN
						next_sreg2<=STATE52;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RD_PTW_PTR_EN_5<='1';
					 ELSE
						next_sreg2<=CRUISEBUFFER_FT;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RD_PTW_PTR_EN_5<='1';
					END IF;
				WHEN CruiseIdle =>
					IF ( CruiseON='1' ) THEN
						next_sreg2<=Cruise_Mode;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RD_PTW_PTR_EN_5<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
					 ELSE
						next_sreg2<=CruiseIdle;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RD_PTW_PTR_EN_5<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
					END IF;
				WHEN FT_HAVE_DATA =>
					next_sreg2<=STATE20;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_RD_PTW_PTR_EN_5<='1';
				WHEN FT_NODATA =>
					next_sreg2<=Cruise_Done_FT;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_RD_PTW_PTR_EN_5<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_CruiseDone<='1';
					next_PTW_CNT_CLR<='1';
				WHEN PINIT_cruise_DLY =>
					next_sreg2<=STATE16;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_RD_PTW_PTR_EN_5<='1';
				WHEN PINT_CALC =>
					IF ( INIT_PED_CALC_DN='1' ) THEN
						next_sreg2<=STATE39;
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_CLR_INIT_PED_CNT<='1';
						next_RD_PTW_PTR_EN_5<='1';
					 ELSE
						next_sreg2<=PINT_CALC;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RD_PTW_PTR_EN_5<='1';
						next_PINIT_CALC_EN<='1';
					END IF;
				WHEN PLOCAL_CALC =>
					IF ( LOC_PED_CALC_DN='1' ) THEN
						next_sreg2<=RestorePTR_FT;
						next_CLR_INIT_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RD_PTW_PTR_EN_5<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RT_PTW_PTR<='1';
						next_CLR_LOC_PED_CNT<='1';
					 ELSE
						next_sreg2<=PLOCAL_CALC;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RD_PTW_PTR_EN_5<='1';
						next_PLOCAL_CALC_EN<='1';
					END IF;
				WHEN RestorePTR_FT =>
					next_sreg2<=STATE18;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RD_PTW_PTR_EN_5<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
				WHEN STATE2 =>
					next_sreg2<=PLOCAL_CALC;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_RD_PTW_PTR_EN_5<='1';
					next_PLOCAL_CALC_EN<='1';
				WHEN STATE14 =>
					next_sreg2<=STATE29;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RD_PTW_PTR_EN_5<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
				WHEN STATE16 =>
					next_sreg2<=PINT_CALC;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_RD_PTW_PTR_EN_5<='1';
					next_PINIT_CALC_EN<='1';
				WHEN STATE17 =>
					next_sreg2<=Cruise_Done_FT;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_RD_PTW_PTR_EN_5<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_CruiseDone<='1';
					next_PTW_CNT_CLR<='1';
				WHEN STATE18 =>
					next_sreg2<=STATE17;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RD_PTW_PTR_EN_5<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
				WHEN STATE20 =>
					next_sreg2<=STATE2;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_RD_PTW_PTR_EN_5<='1';
				WHEN STATE29 =>
					IF ( PTW_DONE='1' ) THEN
						next_sreg2<=FT_NODATA;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RD_PTW_PTR_EN_5<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_NoEventLatch<='1';
					ELSIF ( PTW_DONE='0' ) THEN
						next_sreg2<=STATE14;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RD_PTW_PTR_EN_5<='1';
					END IF;
				WHEN STATE39 =>
					IF ( wait_PG_done='1' ) THEN
						next_sreg2<=STATE40;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RD_PTW_PTR_EN_5<='1';
					 ELSE
						next_sreg2<=STATE39;
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_CLR_INIT_PED_CNT<='1';
						next_RD_PTW_PTR_EN_5<='1';
					END IF;
				WHEN STATE40 =>
					next_sreg2<=STATE67;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_RD_PTW_PTR_EN_5<='1';
				WHEN STATE52 =>
					IF ( WE_DONE='1' ) THEN
						next_sreg2<=STATE14;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RD_PTW_PTR_EN_5<='1';
					ELSIF ( FT_ABOVE_TH='1' AND WE_DONE='0' ) THEN
						next_sreg2<=FT_HAVE_DATA;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RD_PTW_PTR_EN_5<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='1';
						next_SAVE_PTW_PTR_FT<='1';
					ELSIF ( FT_ABOVE_TH='0' AND WE_DONE='0' ) THEN
						next_sreg2<=CRUISEBUFFER_FT;
						next_CLR_INIT_PED_CNT<='0';
						next_CLR_LOC_PED_CNT<='0';
						next_CruiseDone<='0';
						next_NoEventLatch<='0';
						next_PINIT_CALC_EN<='0';
						next_PLOCAL_CALC_EN<='0';
						next_PTW_CNT_CLR<='0';
						next_RT_PTW_PTR<='0';
						next_RT_PTW_PTR_PLOC<='0';
						next_SAVE_PTW_PTR_FT<='0';
						next_RD_PTW_PTR_EN_5<='1';
					END IF;
				WHEN STATE67 =>
					next_sreg2<=CRUISEBUFFER_FT;
					next_CLR_INIT_PED_CNT<='0';
					next_CLR_LOC_PED_CNT<='0';
					next_CruiseDone<='0';
					next_NoEventLatch<='0';
					next_PINIT_CALC_EN<='0';
					next_PLOCAL_CALC_EN<='0';
					next_PTW_CNT_CLR<='0';
					next_RT_PTW_PTR<='0';
					next_RT_PTW_PTR_PLOC<='0';
					next_SAVE_PTW_PTR_FT<='0';
					next_RD_PTW_PTR_EN_5<='1';
				WHEN OTHERS =>
			END CASE;
		END IF;
	END PROCESS;
END BEHAVIOR;

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FT_PROCESSM_CDC_FDC IS
	PORT (MODE : IN std_logic_vector (2 DOWNTO 0);
		CLK,FT_ABOVE_TH,FT_DONE,GO,INIT_PED_CALC_DN,LOC_PED_CALC_DN,NO_EVENT,
			PEAK_WRITE_DONE,PTW_DONE,RESET_N,wait_PG_done,WE_DONE: IN std_logic;
		CLR_INIT_PED_CNT,CLR_LOC_PED_CNT,CLR_PTW_DONE,DEC_PEAK_CNT,FT_GO,
			HOST_BLOCK_INC,IDLE,LatchNoEvenClr,NoEventLatch,NOT_VALID_2,PINIT_CALC_EN,
			PLOCAL_CALC_EN,PR_FIFO_WR_EN,PR_FIFO_WR_EN_TR,PTW_CNT_CLR,RAW_PTW_PTR_EN,
			RD_PTW_PTR_EN_5,RT_PTW_PTR,RT_PTW_PTR_2,RT_PTW_PTR_PLOC,SAVE_PTW_PTR,
			SAVE_PTW_PTR_FT,SEL_CDC_FT_WD_1,SEL_CDC_FT_WD_2,SEL_FDC_AMP_WD_1,
			SEL_FDC_AMP_WD_2,SEL_FDC_SUM_WD_1,SEL_FDC_SUM_WD_2,SEL_RAW_SAMPLE_2,SEL_RS_1,
			SEL_RS_2,SEL_WIN_RAW_WD_1 : OUT std_logic);
END;

ARCHITECTURE BEHAVIOR OF FT_PROCESSM_CDC_FDC IS
	COMPONENT SHELL_FT_PROCESSM_CDC_FDC
		PORT (CLK,FT_ABOVE_TH,FT_DONE,GO,INIT_PED_CALC_DN,LOC_PED_CALC_DN,MODE0,
			MODE1,MODE2,NO_EVENT,PEAK_WRITE_DONE,PTW_DONE,RESET_N,wait_PG_done,WE_DONE: 
			IN std_logic;
			CLR_INIT_PED_CNT,CLR_LOC_PED_CNT,CLR_PTW_DONE,DEC_PEAK_CNT,FT_GO,
				HOST_BLOCK_INC,IDLE,LatchNoEvenClr,NoEventLatch,NOT_VALID_2,PINIT_CALC_EN,
				PLOCAL_CALC_EN,PR_FIFO_WR_EN,PR_FIFO_WR_EN_TR,PTW_CNT_CLR,RAW_PTW_PTR_EN,
				RD_PTW_PTR_EN_5,RT_PTW_PTR,RT_PTW_PTR_2,RT_PTW_PTR_PLOC,SAVE_PTW_PTR,
				SAVE_PTW_PTR_FT,SEL_CDC_FT_WD_1,SEL_CDC_FT_WD_2,SEL_FDC_AMP_WD_1,
				SEL_FDC_AMP_WD_2,SEL_FDC_SUM_WD_1,SEL_FDC_SUM_WD_2,SEL_RAW_SAMPLE_2,SEL_RS_1,
				SEL_RS_2,SEL_WIN_RAW_WD_1 : OUT std_logic);
	END COMPONENT;
BEGIN
	SHELL1_FT_PROCESSM_CDC_FDC : SHELL_FT_PROCESSM_CDC_FDC PORT MAP (CLK=>CLK,
		FT_ABOVE_TH=>FT_ABOVE_TH,FT_DONE=>FT_DONE,GO=>GO,INIT_PED_CALC_DN=>
		INIT_PED_CALC_DN,LOC_PED_CALC_DN=>LOC_PED_CALC_DN,MODE0=>MODE(0),MODE1=>MODE(
		1),MODE2=>MODE(2),NO_EVENT=>NO_EVENT,PEAK_WRITE_DONE=>PEAK_WRITE_DONE,
		PTW_DONE=>PTW_DONE,RESET_N=>RESET_N,wait_PG_done=>wait_PG_done,WE_DONE=>
		WE_DONE,CLR_INIT_PED_CNT=>CLR_INIT_PED_CNT,CLR_LOC_PED_CNT=>CLR_LOC_PED_CNT,
		CLR_PTW_DONE=>CLR_PTW_DONE,DEC_PEAK_CNT=>DEC_PEAK_CNT,FT_GO=>FT_GO,
		HOST_BLOCK_INC=>HOST_BLOCK_INC,IDLE=>IDLE,LatchNoEvenClr=>LatchNoEvenClr,
		NoEventLatch=>NoEventLatch,NOT_VALID_2=>NOT_VALID_2,PINIT_CALC_EN=>
		PINIT_CALC_EN,PLOCAL_CALC_EN=>PLOCAL_CALC_EN,PR_FIFO_WR_EN=>PR_FIFO_WR_EN,
		PR_FIFO_WR_EN_TR=>PR_FIFO_WR_EN_TR,PTW_CNT_CLR=>PTW_CNT_CLR,RAW_PTW_PTR_EN=>
		RAW_PTW_PTR_EN,RD_PTW_PTR_EN_5=>RD_PTW_PTR_EN_5,RT_PTW_PTR=>RT_PTW_PTR,
		RT_PTW_PTR_2=>RT_PTW_PTR_2,RT_PTW_PTR_PLOC=>RT_PTW_PTR_PLOC,SAVE_PTW_PTR=>
		SAVE_PTW_PTR,SAVE_PTW_PTR_FT=>SAVE_PTW_PTR_FT,SEL_CDC_FT_WD_1=>
		SEL_CDC_FT_WD_1,SEL_CDC_FT_WD_2=>SEL_CDC_FT_WD_2,SEL_FDC_AMP_WD_1=>
		SEL_FDC_AMP_WD_1,SEL_FDC_AMP_WD_2=>SEL_FDC_AMP_WD_2,SEL_FDC_SUM_WD_1=>
		SEL_FDC_SUM_WD_1,SEL_FDC_SUM_WD_2=>SEL_FDC_SUM_WD_2,SEL_RAW_SAMPLE_2=>
		SEL_RAW_SAMPLE_2,SEL_RS_1=>SEL_RS_1,SEL_RS_2=>SEL_RS_2,SEL_WIN_RAW_WD_1=>
		SEL_WIN_RAW_WD_1);
END BEHAVIOR;
